magic
tech sky130A
magscale 1 2
timestamp 1640889851
<< obsli1 >>
rect 1104 2159 196943 196945
<< obsm1 >>
rect 14 1980 196955 196976
<< metal2 >>
rect 1490 198656 1546 199456
rect 7378 198656 7434 199456
rect 13266 198656 13322 199456
rect 19338 198656 19394 199456
rect 25226 198656 25282 199456
rect 31114 198656 31170 199456
rect 37002 198656 37058 199456
rect 42890 198656 42946 199456
rect 48962 198656 49018 199456
rect 54850 198656 54906 199456
rect 60738 198656 60794 199456
rect 66626 198656 66682 199456
rect 72698 198656 72754 199456
rect 78586 198656 78642 199456
rect 84474 198656 84530 199456
rect 90362 198656 90418 199456
rect 96434 198656 96490 199456
rect 102322 198656 102378 199456
rect 108210 198656 108266 199456
rect 114098 198656 114154 199456
rect 119986 198656 120042 199456
rect 126058 198656 126114 199456
rect 131946 198656 132002 199456
rect 137834 198656 137890 199456
rect 143722 198656 143778 199456
rect 149794 198656 149850 199456
rect 155682 198656 155738 199456
rect 161570 198656 161626 199456
rect 167458 198656 167514 199456
rect 173530 198656 173586 199456
rect 179418 198656 179474 199456
rect 185306 198656 185362 199456
rect 191194 198656 191250 199456
rect 18 0 74 800
rect 5906 0 5962 800
rect 11794 0 11850 800
rect 17682 0 17738 800
rect 23570 0 23626 800
rect 29642 0 29698 800
rect 35530 0 35586 800
rect 41418 0 41474 800
rect 47306 0 47362 800
rect 53378 0 53434 800
rect 59266 0 59322 800
rect 65154 0 65210 800
rect 71042 0 71098 800
rect 77114 0 77170 800
rect 83002 0 83058 800
rect 88890 0 88946 800
rect 94778 0 94834 800
rect 100666 0 100722 800
rect 106738 0 106794 800
rect 112626 0 112682 800
rect 118514 0 118570 800
rect 124402 0 124458 800
rect 130474 0 130530 800
rect 136362 0 136418 800
rect 142250 0 142306 800
rect 148138 0 148194 800
rect 154210 0 154266 800
rect 160098 0 160154 800
rect 165986 0 166042 800
rect 171874 0 171930 800
rect 177762 0 177818 800
rect 183834 0 183890 800
rect 189722 0 189778 800
rect 195610 0 195666 800
<< obsm2 >>
rect 20 198600 1434 199209
rect 1602 198600 7322 199209
rect 7490 198600 13210 199209
rect 13378 198600 19282 199209
rect 19450 198600 25170 199209
rect 25338 198600 31058 199209
rect 31226 198600 36946 199209
rect 37114 198600 42834 199209
rect 43002 198600 48906 199209
rect 49074 198600 54794 199209
rect 54962 198600 60682 199209
rect 60850 198600 66570 199209
rect 66738 198600 72642 199209
rect 72810 198600 78530 199209
rect 78698 198600 84418 199209
rect 84586 198600 90306 199209
rect 90474 198600 96378 199209
rect 96546 198600 102266 199209
rect 102434 198600 108154 199209
rect 108322 198600 114042 199209
rect 114210 198600 119930 199209
rect 120098 198600 126002 199209
rect 126170 198600 131890 199209
rect 132058 198600 137778 199209
rect 137946 198600 143666 199209
rect 143834 198600 149738 199209
rect 149906 198600 155626 199209
rect 155794 198600 161514 199209
rect 161682 198600 167402 199209
rect 167570 198600 173474 199209
rect 173642 198600 179362 199209
rect 179530 198600 185250 199209
rect 185418 198600 191138 199209
rect 191306 198600 195664 199209
rect 20 856 195664 198600
rect 130 800 5850 856
rect 6018 800 11738 856
rect 11906 800 17626 856
rect 17794 800 23514 856
rect 23682 800 29586 856
rect 29754 800 35474 856
rect 35642 800 41362 856
rect 41530 800 47250 856
rect 47418 800 53322 856
rect 53490 800 59210 856
rect 59378 800 65098 856
rect 65266 800 70986 856
rect 71154 800 77058 856
rect 77226 800 82946 856
rect 83114 800 88834 856
rect 89002 800 94722 856
rect 94890 800 100610 856
rect 100778 800 106682 856
rect 106850 800 112570 856
rect 112738 800 118458 856
rect 118626 800 124346 856
rect 124514 800 130418 856
rect 130586 800 136306 856
rect 136474 800 142194 856
rect 142362 800 148082 856
rect 148250 800 154154 856
rect 154322 800 160042 856
rect 160210 800 165930 856
rect 166098 800 171818 856
rect 171986 800 177706 856
rect 177874 800 183778 856
rect 183946 800 189666 856
rect 189834 800 195554 856
<< metal3 >>
rect 196512 199112 197312 199232
rect 0 192856 800 192976
rect 196512 190408 197312 190528
rect 0 183880 800 184000
rect 196512 181704 197312 181824
rect 0 175176 800 175296
rect 196512 173000 197312 173120
rect 0 166472 800 166592
rect 196512 164296 197312 164416
rect 0 157768 800 157888
rect 196512 155320 197312 155440
rect 0 148792 800 148912
rect 196512 146616 197312 146736
rect 0 140088 800 140208
rect 196512 137912 197312 138032
rect 0 131384 800 131504
rect 196512 129208 197312 129328
rect 0 122680 800 122800
rect 196512 120232 197312 120352
rect 0 113976 800 114096
rect 196512 111528 197312 111648
rect 0 105000 800 105120
rect 196512 102824 197312 102944
rect 0 96296 800 96416
rect 196512 94120 197312 94240
rect 0 87592 800 87712
rect 196512 85144 197312 85264
rect 0 78888 800 79008
rect 196512 76440 197312 76560
rect 0 69912 800 70032
rect 196512 67736 197312 67856
rect 0 61208 800 61328
rect 196512 59032 197312 59152
rect 0 52504 800 52624
rect 196512 50328 197312 50448
rect 0 43800 800 43920
rect 196512 41352 197312 41472
rect 0 34824 800 34944
rect 196512 32648 197312 32768
rect 0 26120 800 26240
rect 196512 23944 197312 24064
rect 0 17416 800 17536
rect 196512 15240 197312 15360
rect 0 8712 800 8832
rect 196512 6264 197312 6384
<< obsm3 >>
rect 800 199032 196432 199205
rect 800 193056 196512 199032
rect 880 192776 196512 193056
rect 800 190608 196512 192776
rect 800 190328 196432 190608
rect 800 184080 196512 190328
rect 880 183800 196512 184080
rect 800 181904 196512 183800
rect 800 181624 196432 181904
rect 800 175376 196512 181624
rect 880 175096 196512 175376
rect 800 173200 196512 175096
rect 800 172920 196432 173200
rect 800 166672 196512 172920
rect 880 166392 196512 166672
rect 800 164496 196512 166392
rect 800 164216 196432 164496
rect 800 157968 196512 164216
rect 880 157688 196512 157968
rect 800 155520 196512 157688
rect 800 155240 196432 155520
rect 800 148992 196512 155240
rect 880 148712 196512 148992
rect 800 146816 196512 148712
rect 800 146536 196432 146816
rect 800 140288 196512 146536
rect 880 140008 196512 140288
rect 800 138112 196512 140008
rect 800 137832 196432 138112
rect 800 131584 196512 137832
rect 880 131304 196512 131584
rect 800 129408 196512 131304
rect 800 129128 196432 129408
rect 800 122880 196512 129128
rect 880 122600 196512 122880
rect 800 120432 196512 122600
rect 800 120152 196432 120432
rect 800 114176 196512 120152
rect 880 113896 196512 114176
rect 800 111728 196512 113896
rect 800 111448 196432 111728
rect 800 105200 196512 111448
rect 880 104920 196512 105200
rect 800 103024 196512 104920
rect 800 102744 196432 103024
rect 800 96496 196512 102744
rect 880 96216 196512 96496
rect 800 94320 196512 96216
rect 800 94040 196432 94320
rect 800 87792 196512 94040
rect 880 87512 196512 87792
rect 800 85344 196512 87512
rect 800 85064 196432 85344
rect 800 79088 196512 85064
rect 880 78808 196512 79088
rect 800 76640 196512 78808
rect 800 76360 196432 76640
rect 800 70112 196512 76360
rect 880 69832 196512 70112
rect 800 67936 196512 69832
rect 800 67656 196432 67936
rect 800 61408 196512 67656
rect 880 61128 196512 61408
rect 800 59232 196512 61128
rect 800 58952 196432 59232
rect 800 52704 196512 58952
rect 880 52424 196512 52704
rect 800 50528 196512 52424
rect 800 50248 196432 50528
rect 800 44000 196512 50248
rect 880 43720 196512 44000
rect 800 41552 196512 43720
rect 800 41272 196432 41552
rect 800 35024 196512 41272
rect 880 34744 196512 35024
rect 800 32848 196512 34744
rect 800 32568 196432 32848
rect 800 26320 196512 32568
rect 880 26040 196512 26320
rect 800 24144 196512 26040
rect 800 23864 196432 24144
rect 800 17616 196512 23864
rect 880 17336 196512 17616
rect 800 15440 196512 17336
rect 800 15160 196432 15440
rect 800 8912 196512 15160
rect 880 8632 196512 8912
rect 800 6464 196512 8632
rect 800 6184 196432 6464
rect 800 1939 196512 6184
<< metal4 >>
rect 4208 2128 4528 196976
rect 19568 2128 19888 196976
rect 34928 2128 35248 196976
rect 50288 2128 50608 196976
rect 65648 2128 65968 196976
rect 81008 2128 81328 196976
rect 96368 2128 96688 196976
rect 111728 2128 112048 196976
rect 127088 2128 127408 196976
rect 142448 2128 142768 196976
rect 157808 2128 158128 196976
rect 173168 2128 173488 196976
rect 188528 2128 188848 196976
<< obsm4 >>
rect 34651 2048 34848 179893
rect 35328 2048 50208 179893
rect 50688 2048 65568 179893
rect 66048 2048 80928 179893
rect 81408 2048 96288 179893
rect 96768 2048 111648 179893
rect 112128 2048 127008 179893
rect 127488 2048 142368 179893
rect 142848 2048 157728 179893
rect 158208 2048 167565 179893
rect 34651 1939 167565 2048
<< labels >>
rlabel metal3 s 196512 50328 197312 50448 6 io_oeb
port 1 nsew signal output
rlabel metal2 s 90362 198656 90418 199456 6 io_out
port 2 nsew signal output
rlabel metal3 s 0 78888 800 79008 6 irq[0]
port 3 nsew signal output
rlabel metal2 s 131946 198656 132002 199456 6 irq[1]
port 4 nsew signal output
rlabel metal2 s 1490 198656 1546 199456 6 irq[2]
port 5 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 la_data_in
port 6 nsew signal input
rlabel metal4 s 4208 2128 4528 196976 6 vccd1
port 7 nsew power input
rlabel metal4 s 34928 2128 35248 196976 6 vccd1
port 7 nsew power input
rlabel metal4 s 65648 2128 65968 196976 6 vccd1
port 7 nsew power input
rlabel metal4 s 96368 2128 96688 196976 6 vccd1
port 7 nsew power input
rlabel metal4 s 127088 2128 127408 196976 6 vccd1
port 7 nsew power input
rlabel metal4 s 157808 2128 158128 196976 6 vccd1
port 7 nsew power input
rlabel metal4 s 188528 2128 188848 196976 6 vccd1
port 7 nsew power input
rlabel metal4 s 19568 2128 19888 196976 6 vssd1
port 8 nsew ground input
rlabel metal4 s 50288 2128 50608 196976 6 vssd1
port 8 nsew ground input
rlabel metal4 s 81008 2128 81328 196976 6 vssd1
port 8 nsew ground input
rlabel metal4 s 111728 2128 112048 196976 6 vssd1
port 8 nsew ground input
rlabel metal4 s 142448 2128 142768 196976 6 vssd1
port 8 nsew ground input
rlabel metal4 s 173168 2128 173488 196976 6 vssd1
port 8 nsew ground input
rlabel metal3 s 0 157768 800 157888 6 wb_clk_i
port 9 nsew signal input
rlabel metal3 s 0 105000 800 105120 6 wb_rst_i
port 10 nsew signal input
rlabel metal2 s 84474 198656 84530 199456 6 wbs_ack_o
port 11 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 wbs_adr_i[0]
port 12 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 wbs_adr_i[10]
port 13 nsew signal input
rlabel metal2 s 179418 198656 179474 199456 6 wbs_adr_i[11]
port 14 nsew signal input
rlabel metal2 s 160098 0 160154 800 6 wbs_adr_i[12]
port 15 nsew signal input
rlabel metal3 s 196512 173000 197312 173120 6 wbs_adr_i[13]
port 16 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 wbs_adr_i[14]
port 17 nsew signal input
rlabel metal2 s 177762 0 177818 800 6 wbs_adr_i[15]
port 18 nsew signal input
rlabel metal3 s 196512 155320 197312 155440 6 wbs_adr_i[16]
port 19 nsew signal input
rlabel metal2 s 114098 198656 114154 199456 6 wbs_adr_i[17]
port 20 nsew signal input
rlabel metal2 s 54850 198656 54906 199456 6 wbs_adr_i[18]
port 21 nsew signal input
rlabel metal3 s 196512 181704 197312 181824 6 wbs_adr_i[19]
port 22 nsew signal input
rlabel metal2 s 72698 198656 72754 199456 6 wbs_adr_i[1]
port 23 nsew signal input
rlabel metal3 s 0 148792 800 148912 6 wbs_adr_i[20]
port 24 nsew signal input
rlabel metal2 s 154210 0 154266 800 6 wbs_adr_i[21]
port 25 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 wbs_adr_i[22]
port 26 nsew signal input
rlabel metal2 s 119986 198656 120042 199456 6 wbs_adr_i[23]
port 27 nsew signal input
rlabel metal2 s 136362 0 136418 800 6 wbs_adr_i[24]
port 28 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_adr_i[25]
port 29 nsew signal input
rlabel metal2 s 102322 198656 102378 199456 6 wbs_adr_i[26]
port 30 nsew signal input
rlabel metal3 s 196512 15240 197312 15360 6 wbs_adr_i[27]
port 31 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 wbs_adr_i[28]
port 32 nsew signal input
rlabel metal2 s 25226 198656 25282 199456 6 wbs_adr_i[29]
port 33 nsew signal input
rlabel metal3 s 0 175176 800 175296 6 wbs_adr_i[2]
port 34 nsew signal input
rlabel metal2 s 167458 198656 167514 199456 6 wbs_adr_i[30]
port 35 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 wbs_adr_i[31]
port 36 nsew signal input
rlabel metal3 s 196512 23944 197312 24064 6 wbs_adr_i[3]
port 37 nsew signal input
rlabel metal3 s 196512 164296 197312 164416 6 wbs_adr_i[4]
port 38 nsew signal input
rlabel metal3 s 196512 137912 197312 138032 6 wbs_adr_i[5]
port 39 nsew signal input
rlabel metal3 s 196512 120232 197312 120352 6 wbs_adr_i[6]
port 40 nsew signal input
rlabel metal3 s 196512 111528 197312 111648 6 wbs_adr_i[7]
port 41 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 wbs_adr_i[8]
port 42 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 wbs_adr_i[9]
port 43 nsew signal input
rlabel metal3 s 196512 190408 197312 190528 6 wbs_cyc_i
port 44 nsew signal input
rlabel metal3 s 0 166472 800 166592 6 wbs_dat_i[0]
port 45 nsew signal input
rlabel metal2 s 108210 198656 108266 199456 6 wbs_dat_i[10]
port 46 nsew signal input
rlabel metal3 s 196512 76440 197312 76560 6 wbs_dat_i[11]
port 47 nsew signal input
rlabel metal3 s 196512 85144 197312 85264 6 wbs_dat_i[12]
port 48 nsew signal input
rlabel metal2 s 78586 198656 78642 199456 6 wbs_dat_i[13]
port 49 nsew signal input
rlabel metal2 s 126058 198656 126114 199456 6 wbs_dat_i[14]
port 50 nsew signal input
rlabel metal2 s 185306 198656 185362 199456 6 wbs_dat_i[15]
port 51 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 wbs_dat_i[16]
port 52 nsew signal input
rlabel metal3 s 196512 6264 197312 6384 6 wbs_dat_i[17]
port 53 nsew signal input
rlabel metal2 s 183834 0 183890 800 6 wbs_dat_i[18]
port 54 nsew signal input
rlabel metal3 s 0 122680 800 122800 6 wbs_dat_i[19]
port 55 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_dat_i[1]
port 56 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 wbs_dat_i[20]
port 57 nsew signal input
rlabel metal2 s 195610 0 195666 800 6 wbs_dat_i[21]
port 58 nsew signal input
rlabel metal3 s 196512 199112 197312 199232 6 wbs_dat_i[22]
port 59 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 wbs_dat_i[23]
port 60 nsew signal input
rlabel metal2 s 130474 0 130530 800 6 wbs_dat_i[24]
port 61 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 wbs_dat_i[25]
port 62 nsew signal input
rlabel metal3 s 196512 32648 197312 32768 6 wbs_dat_i[26]
port 63 nsew signal input
rlabel metal2 s 66626 198656 66682 199456 6 wbs_dat_i[27]
port 64 nsew signal input
rlabel metal3 s 0 192856 800 192976 6 wbs_dat_i[28]
port 65 nsew signal input
rlabel metal2 s 171874 0 171930 800 6 wbs_dat_i[29]
port 66 nsew signal input
rlabel metal2 s 19338 198656 19394 199456 6 wbs_dat_i[2]
port 67 nsew signal input
rlabel metal3 s 0 43800 800 43920 6 wbs_dat_i[30]
port 68 nsew signal input
rlabel metal2 s 143722 198656 143778 199456 6 wbs_dat_i[31]
port 69 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 wbs_dat_i[3]
port 70 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_i[4]
port 71 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 wbs_dat_i[5]
port 72 nsew signal input
rlabel metal2 s 165986 0 166042 800 6 wbs_dat_i[6]
port 73 nsew signal input
rlabel metal3 s 196512 94120 197312 94240 6 wbs_dat_i[7]
port 74 nsew signal input
rlabel metal3 s 196512 41352 197312 41472 6 wbs_dat_i[8]
port 75 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 wbs_dat_i[9]
port 76 nsew signal input
rlabel metal3 s 0 183880 800 184000 6 wbs_dat_o[0]
port 77 nsew signal output
rlabel metal3 s 0 140088 800 140208 6 wbs_dat_o[10]
port 78 nsew signal output
rlabel metal3 s 0 131384 800 131504 6 wbs_dat_o[11]
port 79 nsew signal output
rlabel metal3 s 196512 59032 197312 59152 6 wbs_dat_o[12]
port 80 nsew signal output
rlabel metal3 s 196512 129208 197312 129328 6 wbs_dat_o[13]
port 81 nsew signal output
rlabel metal2 s 142250 0 142306 800 6 wbs_dat_o[14]
port 82 nsew signal output
rlabel metal3 s 196512 146616 197312 146736 6 wbs_dat_o[15]
port 83 nsew signal output
rlabel metal3 s 0 52504 800 52624 6 wbs_dat_o[16]
port 84 nsew signal output
rlabel metal2 s 42890 198656 42946 199456 6 wbs_dat_o[17]
port 85 nsew signal output
rlabel metal3 s 0 96296 800 96416 6 wbs_dat_o[18]
port 86 nsew signal output
rlabel metal2 s 18 0 74 800 6 wbs_dat_o[19]
port 87 nsew signal output
rlabel metal2 s 106738 0 106794 800 6 wbs_dat_o[1]
port 88 nsew signal output
rlabel metal2 s 48962 198656 49018 199456 6 wbs_dat_o[20]
port 89 nsew signal output
rlabel metal2 s 96434 198656 96490 199456 6 wbs_dat_o[21]
port 90 nsew signal output
rlabel metal2 s 149794 198656 149850 199456 6 wbs_dat_o[22]
port 91 nsew signal output
rlabel metal2 s 13266 198656 13322 199456 6 wbs_dat_o[23]
port 92 nsew signal output
rlabel metal3 s 0 113976 800 114096 6 wbs_dat_o[24]
port 93 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[25]
port 94 nsew signal output
rlabel metal2 s 173530 198656 173586 199456 6 wbs_dat_o[26]
port 95 nsew signal output
rlabel metal2 s 137834 198656 137890 199456 6 wbs_dat_o[27]
port 96 nsew signal output
rlabel metal2 s 77114 0 77170 800 6 wbs_dat_o[28]
port 97 nsew signal output
rlabel metal2 s 191194 198656 191250 199456 6 wbs_dat_o[29]
port 98 nsew signal output
rlabel metal2 s 189722 0 189778 800 6 wbs_dat_o[2]
port 99 nsew signal output
rlabel metal2 s 31114 198656 31170 199456 6 wbs_dat_o[30]
port 100 nsew signal output
rlabel metal3 s 0 87592 800 87712 6 wbs_dat_o[31]
port 101 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 wbs_dat_o[3]
port 102 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 wbs_dat_o[4]
port 103 nsew signal output
rlabel metal2 s 88890 0 88946 800 6 wbs_dat_o[5]
port 104 nsew signal output
rlabel metal3 s 196512 102824 197312 102944 6 wbs_dat_o[6]
port 105 nsew signal output
rlabel metal2 s 94778 0 94834 800 6 wbs_dat_o[7]
port 106 nsew signal output
rlabel metal2 s 161570 198656 161626 199456 6 wbs_dat_o[8]
port 107 nsew signal output
rlabel metal2 s 155682 198656 155738 199456 6 wbs_dat_o[9]
port 108 nsew signal output
rlabel metal2 s 37002 198656 37058 199456 6 wbs_sel_i[0]
port 109 nsew signal input
rlabel metal2 s 60738 198656 60794 199456 6 wbs_sel_i[1]
port 110 nsew signal input
rlabel metal2 s 112626 0 112682 800 6 wbs_sel_i[2]
port 111 nsew signal input
rlabel metal3 s 0 69912 800 70032 6 wbs_sel_i[3]
port 112 nsew signal input
rlabel metal2 s 7378 198656 7434 199456 6 wbs_stb_i
port 113 nsew signal input
rlabel metal3 s 196512 67736 197312 67856 6 wbs_we_i
port 114 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 197312 199456
string LEFview TRUE
string GDS_FILE /project/sky130-openlane/runs/subservient_wrapped/results/magic/subservient_wrapped.gds
string GDS_END 83861520
string GDS_START 772160
<< end >>

